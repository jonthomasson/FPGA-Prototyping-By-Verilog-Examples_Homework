library verilog;
use verilog.vl_types.all;
entity bin_counter_tb is
end bin_counter_tb;
