library verilog;
use verilog.vl_types.all;
entity occupancy_counter_tb is
end occupancy_counter_tb;
