library verilog;
use verilog.vl_types.all;
entity square_wave_tb is
end square_wave_tb;
