// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module font_rom
   (
    input wire clk,
    input wire [14:0] addr,
    output reg [7:0] data
   );
   
   // signal declaration
   reg [14:0] addr_reg; 

   // body
   always @(posedge clk) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)
         //code x00
         15'h0000: data = 8'b00000000; // 
         15'h0001: data = 8'b00000000; // 
         15'h0002: data = 8'b00000000; // 
         15'h0003: data = 8'b00000000; // 
         15'h0004: data = 8'b00000000; // 
         15'h0005: data = 8'b00000000; // 
         15'h0006: data = 8'b00000000; // 
         15'h0007: data = 8'b00000000; // 
         15'h0008: data = 8'b00000000; // 
         15'h0009: data = 8'b00000000; // 
         15'h000a: data = 8'b00000000; // 
         15'h000b: data = 8'b00000000; // 
         15'h000c: data = 8'b00000000; // 
         15'h000d: data = 8'b00000000; // 
         15'h000e: data = 8'b00000000; // 
         15'h000f: data = 8'b00000000; // 
         15'h0010: data = 8'b00000000; // 
         15'h0011: data = 8'b00000000; // 
         15'h0012: data = 8'b00000000; //  
         15'h0013: data = 8'b00000000; // 
         15'h0014: data = 8'b00000000; // 
         15'h0015: data = 8'b00000000; //
         15'h0016: data = 8'b00000000; // 
         15'h0017: data = 8'b00000000; // 
         15'h0018: data = 8'b00000000; // 
         15'h0019: data = 8'b00000000; // 
         15'h001a: data = 8'b00000000; // 
         15'h001b: data = 8'b00000000; // 
         15'h001c: data = 8'b00000000; // 
         15'h001d: data = 8'b00000000; // 
         15'h001e: data = 8'b00000000; // 
         15'h001f: data = 8'b00000000; // 
         15'h0020: data = 8'b00000000; // 
         15'h0021: data = 8'b00000000; // 
         15'h0022: data = 8'b00000000; //  
         15'h0023: data = 8'b00000000; // 
         15'h0024: data = 8'b00000000; // 
         15'h0025: data = 8'b00000000; // 
         15'h0026: data = 8'b00000000; // 
         15'h0027: data = 8'b00000000; // 
         15'h0028: data = 8'b00000000; // 
         15'h0029: data = 8'b00000000; // 
         15'h002a: data = 8'b00000000; // 
         15'h002b: data = 8'b00000000; //  
         15'h002c: data = 8'b00000000; // 
         15'h002d: data = 8'b00000000; // 
         15'h002e: data = 8'b00000000; // 
         15'h002f: data = 8'b00000000; // 
         15'h0030: data = 8'b00000000; // 
         15'h0031: data = 8'b00000000; // 
         15'h0032: data = 8'b00000000; // 
         15'h0033: data = 8'b00000000; // 
         15'h0034: data = 8'b00000000; //  
         15'h0035: data = 8'b00000000; // 
         15'h0036: data = 8'b00000000; // 
         15'h0037: data = 8'b00000000; // 
         15'h0038: data = 8'b00000000; // 
         15'h0039: data = 8'b00000000; //  
         15'h003a: data = 8'b11111111; // ********  
         15'h003b: data = 8'b11111111; // ********
         15'h003c: data = 8'b00000000; // 
         15'h003d: data = 8'b00000000; // 
         15'h003e: data = 8'b00000000; // 
         15'h003f: data = 8'b00000000; // 
         //code x01
         15'h0100: data = 8'b00000000; // 
         15'h0101: data = 8'b00000000; // 
         15'h0102: data = 8'b00011111; //    *****
         15'h0103: data = 8'b00011111; //    *****
         15'h0104: data = 8'b00011000; //    **
         15'h0105: data = 8'b00011000; //    **
         15'h0106: data = 8'b00011000; //    **
         15'h0107: data = 8'b00011000; //    **
         15'h0108: data = 8'b00011000; //    **
         15'h0109: data = 8'b00011000; //    **
         15'h010a: data = 8'b00011000; //    **
         15'h010b: data = 8'b00011000; //    **
         15'h010c: data = 8'b00011000; //    **
         15'h010d: data = 8'b00011000; //    **
         15'h010e: data = 8'b00011000; //    **
         15'h010f: data = 8'b00011000; //    **
         15'h0110: data = 8'b00011000; //    **
         15'h0111: data = 8'b00011000; //    **
         15'h0112: data = 8'b00011000; //    **
         15'h0113: data = 8'b00011000; //    **
         15'h0114: data = 8'b00011000; //    **
         15'h0115: data = 8'b00011000; //    **
         15'h0116: data = 8'b00011000; //    **
         15'h0117: data = 8'b00011000; //    **
         15'h0118: data = 8'b00011000; //    **
         15'h0119: data = 8'b00011000; //    **
         15'h011a: data = 8'b00011000; //    **
         15'h011b: data = 8'b00011000; //    **
         15'h011c: data = 8'b00011000; //    **
         15'h011d: data = 8'b00011000; //    **
         15'h011e: data = 8'b00011000; //    **
         15'h011f: data = 8'b00011000; //    **
         15'h0120: data = 8'b00011000; //    **
         15'h0121: data = 8'b00011000; //    **
         15'h0122: data = 8'b00011000; //    **
         15'h0123: data = 8'b00011000; //    **
         15'h0124: data = 8'b00011000; //    **
         15'h0125: data = 8'b00011000; //    **
         15'h0126: data = 8'b00011000; //    **
         15'h0127: data = 8'b00011000; //    **
         15'h0128: data = 8'b00011000; //    **
         15'h0129: data = 8'b00011000; //    **
         15'h012a: data = 8'b00011000; //    **
         15'h012b: data = 8'b00011000; //    **
         15'h012c: data = 8'b00011000; //    **
         15'h012d: data = 8'b00011000; //    **
         15'h012e: data = 8'b00011000; //    **
         15'h012f: data = 8'b00011000; //    **
         15'h0130: data = 8'b00011000; //    **
         15'h0131: data = 8'b00011000; //    **
         15'h0132: data = 8'b00011000; //    **
         15'h0133: data = 8'b00011000; //    **
         15'h0134: data = 8'b00011000; //    **
         15'h0135: data = 8'b00011000; //    **
         15'h0136: data = 8'b00011000; //    **
         15'h0137: data = 8'b00011000; //    **
         15'h0138: data = 8'b00011000; //    **
         15'h0139: data = 8'b00011000; //    **
         15'h013a: data = 8'b11111000; // *****  
         15'h013b: data = 8'b11111000; // *****
         15'h013c: data = 8'b00000000; // 
         15'h013d: data = 8'b00000000; // 
         15'h013e: data = 8'b00000000; // 
         15'h013f: data = 8'b00000000; // 
         //code x10
         15'h1000: data = 8'b00000000; // 
         15'h1001: data = 8'b00000000; // 
         15'h1002: data = 8'b11111000; // *****
         15'h1003: data = 8'b11111000; // *****
         15'h1004: data = 8'b00011000; //    **
         15'h1005: data = 8'b00011000; //    **
         15'h1006: data = 8'b00011000; //    **
         15'h1007: data = 8'b00011000; //    **
         15'h1008: data = 8'b00011000; //    **
         15'h1009: data = 8'b00011000; //    **
         15'h100a: data = 8'b00011000; //    **
         15'h100b: data = 8'b00011000; //    **
         15'h100c: data = 8'b00011000; //    **
         15'h100d: data = 8'b00011000; //    **
         15'h100e: data = 8'b00011000; //    **
         15'h100f: data = 8'b00011000; //    **
         15'h1010: data = 8'b00011000; //    **
         15'h1011: data = 8'b00011000; //    **
         15'h1012: data = 8'b00011000; //    **
         15'h1013: data = 8'b00011000; //    **
         15'h1014: data = 8'b00011000; //    **
         15'h1015: data = 8'b00011000; //    **
         15'h1016: data = 8'b00011000; //    **
         15'h1017: data = 8'b00011000; //    **
         15'h1018: data = 8'b00011000; //    **
         15'h1019: data = 8'b00011000; //    **
         15'h101a: data = 8'b00011000; //    **
         15'h101b: data = 8'b00011000; //    **
         15'h101c: data = 8'b00011000; //    **
         15'h101d: data = 8'b00011000; //    **
         15'h101e: data = 8'b00011000; //    **
         15'h101f: data = 8'b00011000; //    **
         15'h1020: data = 8'b00011000; //    **
         15'h1021: data = 8'b00011000; //    **
         15'h1022: data = 8'b00011000; //    **
         15'h1023: data = 8'b00011000; //    **
         15'h1024: data = 8'b00011000; //    **
         15'h1025: data = 8'b00011000; //    **
         15'h1026: data = 8'b00011000; //    **
         15'h1027: data = 8'b00011000; //    **
         15'h1028: data = 8'b00011000; //    **
         15'h1029: data = 8'b00011000; //    **
         15'h102a: data = 8'b00011000; //    **
         15'h102b: data = 8'b00011000; //    **
         15'h102c: data = 8'b00011000; //    **
         15'h102d: data = 8'b00011000; //    **
         15'h102e: data = 8'b00011000; //    **
         15'h102f: data = 8'b00011000; //    **
         15'h1030: data = 8'b00011000; //    **
         15'h1031: data = 8'b00011000; //    **
         15'h1032: data = 8'b00011000; //    **
         15'h1033: data = 8'b00011000; //    **
         15'h1034: data = 8'b00011000; //    **
         15'h1035: data = 8'b00011000; //    **
         15'h1036: data = 8'b00011000; //    **
         15'h1037: data = 8'b00011000; //    **
         15'h1038: data = 8'b00011000; //    **
         15'h1039: data = 8'b00011000; //    **
         15'h103a: data = 8'b00011111; //    *****  
         15'h103b: data = 8'b00011111; //    *****
         15'h103c: data = 8'b00000000; // 
         15'h103d: data = 8'b00000000; // 
         15'h103e: data = 8'b00000000; // 
         15'h103f: data = 8'b00000000; // 
         //code x11
         15'h1100: data = 8'b00000000; // 
         15'h1101: data = 8'b00000000; // 
         15'h1102: data = 8'b11111111; // ********
         15'h1103: data = 8'b11111111; // ********
         15'h1104: data = 8'b00000000; // 
         15'h1105: data = 8'b00000000; // 
         15'h1106: data = 8'b00000000; // 
         15'h1107: data = 8'b00000000; // 
         15'h1108: data = 8'b00000000; // 
         15'h1109: data = 8'b00000000; // 
         15'h110a: data = 8'b00000000; // 
         15'h110b: data = 8'b00000000; // 
         15'h110c: data = 8'b00000000; // 
         15'h110d: data = 8'b00000000; // 
         15'h110e: data = 8'b00000000; // 
         15'h110f: data = 8'b00000000; // 
         15'h1110: data = 8'b00000000; // 
         15'h1111: data = 8'b00000000; // 
         15'h1112: data = 8'b00000000; //  
         15'h1113: data = 8'b00000000; // 
         15'h1114: data = 8'b00000000; // 
         15'h1115: data = 8'b00000000; //
         15'h1116: data = 8'b00000000; // 
         15'h1117: data = 8'b00000000; // 
         15'h1118: data = 8'b00000000; // 
         15'h1119: data = 8'b00000000; // 
         15'h111a: data = 8'b00000000; // 
         15'h111b: data = 8'b00000000; // 
         15'h111c: data = 8'b00000000; // 
         15'h111d: data = 8'b00000000; // 
         15'h111e: data = 8'b00000000; // 
         15'h111f: data = 8'b00000000; // 
         15'h1120: data = 8'b00000000; // 
         15'h1121: data = 8'b00000000; // 
         15'h1122: data = 8'b00000000; //  
         15'h1123: data = 8'b00000000; // 
         15'h1124: data = 8'b00000000; // 
         15'h1125: data = 8'b00000000; // 
         15'h1126: data = 8'b00000000; // 
         15'h1127: data = 8'b00000000; // 
         15'h1128: data = 8'b00000000; // 
         15'h1129: data = 8'b00000000; // 
         15'h112a: data = 8'b00000000; // 
         15'h112b: data = 8'b00000000; //  
         15'h112c: data = 8'b00000000; // 
         15'h112d: data = 8'b00000000; // 
         15'h112e: data = 8'b00000000; // 
         15'h112f: data = 8'b00000000; // 
         15'h1130: data = 8'b00000000; // 
         15'h1131: data = 8'b00000000; // 
         15'h1132: data = 8'b00000000; // 
         15'h1133: data = 8'b00000000; // 
         15'h1134: data = 8'b00000000; //  
         15'h1135: data = 8'b00000000; // 
         15'h1136: data = 8'b00000000; // 
         15'h1137: data = 8'b00000000; // 
         15'h1138: data = 8'b00000000; // 
         15'h1139: data = 8'b00000000; //  
         15'h113a: data = 8'b00000000; //  
         15'h113b: data = 8'b00000000; // 
         15'h113c: data = 8'b00000000; // 
         15'h113d: data = 8'b00000000; // 
         15'h113e: data = 8'b00000000; // 
         15'h113f: data = 8'b00000000; // 
   endcase  
   	       
endmodule      
