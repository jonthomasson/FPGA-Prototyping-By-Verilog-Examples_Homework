library verilog;
use verilog.vl_types.all;
entity bcd2bin_tb is
end bcd2bin_tb;
