library verilog;
use verilog.vl_types.all;
entity shiftregister_test is
end shiftregister_test;
