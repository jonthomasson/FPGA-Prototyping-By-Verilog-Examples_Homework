library verilog;
use verilog.vl_types.all;
entity edge_detect_moore_tb is
end edge_detect_moore_tb;
